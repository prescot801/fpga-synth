module note2dds(CLK, NOTE, ADDER);

input wire CLK;
input wire [6:0] NOTE;
output reg [31:0] ADDER;

initial begin
	ADDER = 32'd0;
end

always @ (posedge CLK) begin
	case(NOTE)
		7'd000: ADDER <= 32'd0702;
		7'd001: ADDER <= 32'd0702;
		7'd002: ADDER <= 32'd0702;
		7'd003: ADDER <= 32'd0702;
		7'd004: ADDER <= 32'd0702;
		7'd005: ADDER <= 32'd0702;
		7'd006: ADDER <= 32'd0702;
		7'd007: ADDER <= 32'd0702;
		7'd008: ADDER <= 32'd0702;
		7'd009: ADDER <= 32'd0702;
		7'd010: ADDER <= 32'd0702;
		7'd011: ADDER <= 32'd0702;
		7'd012: ADDER <= 32'd0702;
		7'd013: ADDER <= 32'd0744;
		7'd014: ADDER <= 32'd0788;
		7'd015: ADDER <= 32'd0835;
		7'd016: ADDER <= 32'd0885;
		7'd017: ADDER <= 32'd0937;
		7'd018: ADDER <= 32'd0993;
		7'd019: ADDER <= 32'd01052;
		7'd020: ADDER <= 32'd01115;
		7'd021: ADDER <= 32'd01181;
		7'd022: ADDER <= 32'd01251;
		7'd023: ADDER <= 32'd01326;
		7'd024: ADDER <= 32'd01405;
		7'd025: ADDER <= 32'd01488;
		7'd026: ADDER <= 32'd01577;
		7'd027: ADDER <= 32'd01670;
		7'd028: ADDER <= 32'd01770;
		7'd029: ADDER <= 32'd01875;
		7'd030: ADDER <= 32'd01986;
		7'd031: ADDER <= 32'd02105;
		7'd032: ADDER <= 32'd02230;
		7'd033: ADDER <= 32'd02362;
		7'd034: ADDER <= 32'd02503;
		7'd035: ADDER <= 32'd02652;
		7'd036: ADDER <= 32'd02809;
		7'd037: ADDER <= 32'd02976;
		7'd038: ADDER <= 32'd03153;
		7'd039: ADDER <= 32'd03341;
		7'd040: ADDER <= 32'd03539;
		7'd041: ADDER <= 32'd03750;
		7'd042: ADDER <= 32'd03973;
		7'd043: ADDER <= 32'd04209;
		7'd044: ADDER <= 32'd04459;
		7'd045: ADDER <= 32'd04724;
		7'd046: ADDER <= 32'd05005;
		7'd047: ADDER <= 32'd05303;
		7'd048: ADDER <= 32'd05618;
		7'd049: ADDER <= 32'd05952;
		7'd050: ADDER <= 32'd06306;
		7'd051: ADDER <= 32'd06681;
		7'd052: ADDER <= 32'd07079;
		7'd053: ADDER <= 32'd07500;
		7'd054: ADDER <= 32'd07946;
		7'd055: ADDER <= 32'd08418;
		7'd056: ADDER <= 32'd08919;
		7'd057: ADDER <= 32'd09449;
		7'd058: ADDER <= 32'd010011;
		7'd059: ADDER <= 32'd010606;
		7'd060: ADDER <= 32'd011237;
		7'd061: ADDER <= 32'd011905;
		7'd062: ADDER <= 32'd012613;
		7'd063: ADDER <= 32'd013363;
		7'd064: ADDER <= 32'd014157;
		7'd065: ADDER <= 32'd014999;
		7'd066: ADDER <= 32'd015891;
		7'd067: ADDER <= 32'd016836;
		7'd068: ADDER <= 32'd017837;
		7'd069: ADDER <= 32'd018898;
		7'd070: ADDER <= 32'd020022;
		7'd071: ADDER <= 32'd021212;
		7'd072: ADDER <= 32'd022473;
		7'd073: ADDER <= 32'd023810;
		7'd074: ADDER <= 32'd025226;
		7'd075: ADDER <= 32'd026726;
		7'd076: ADDER <= 32'd028315;
		7'd077: ADDER <= 32'd029998;
		7'd078: ADDER <= 32'd031782;
		7'd079: ADDER <= 32'd033672;
		7'd080: ADDER <= 32'd035674;
		7'd081: ADDER <= 32'd037796;
		7'd082: ADDER <= 32'd040043;
		7'd083: ADDER <= 32'd042424;
		7'd084: ADDER <= 32'd044947;
		7'd085: ADDER <= 32'd047620;
		7'd086: ADDER <= 32'd050451;
		7'd087: ADDER <= 32'd053451;
		7'd088: ADDER <= 32'd056630;
		7'd089: ADDER <= 32'd059997;
		7'd090: ADDER <= 32'd063565;
		7'd091: ADDER <= 32'd067344;
		7'd092: ADDER <= 32'd071349;
		7'd093: ADDER <= 32'd075591;
		7'd094: ADDER <= 32'd080086;
		7'd095: ADDER <= 32'd084849;
		7'd096: ADDER <= 32'd089894;
		7'd097: ADDER <= 32'd095239;
		7'd098: ADDER <= 32'd0100902;
		7'd099: ADDER <= 32'd0106902;
		7'd0100: ADDER <= 32'd0113259;
		7'd0101: ADDER <= 32'd0119994;
		7'd0102: ADDER <= 32'd0127129;
		7'd0103: ADDER <= 32'd0134689;
		7'd0104: ADDER <= 32'd0142698;
		7'd0105: ADDER <= 32'd0151183;
		7'd0106: ADDER <= 32'd0160173;
		7'd0107: ADDER <= 32'd0169697;
		7'd0108: ADDER <= 32'd0179788;
		7'd0109: ADDER <= 32'd0190478;
		7'd0110: ADDER <= 32'd0201805;
		7'd0111: ADDER <= 32'd0213805;
		7'd0112: ADDER <= 32'd0226518;
		7'd0113: ADDER <= 32'd0239988;
		7'd0114: ADDER <= 32'd0254258;
		7'd0115: ADDER <= 32'd0269377;
		7'd0116: ADDER <= 32'd0285395;
		7'd0117: ADDER <= 32'd0302366;
		7'd0118: ADDER <= 32'd0320345;
		7'd0119: ADDER <= 32'd0339394;
		7'd0120: ADDER <= 32'd0359575;
		7'd0121: ADDER <= 32'd0380957;
		7'd0122: ADDER <= 32'd0403610;
		7'd0123: ADDER <= 32'd0427610;
		7'd0124: ADDER <= 32'd0453037;
		7'd0125: ADDER <= 32'd0479976;
		7'd0126: ADDER <= 32'd0508516;
		7'd0127: ADDER <= 32'd0538754;
	endcase
end

endmodule

module lin2exp_t(in_data, out_data);

input wire [6:0] in_data;
output wire [31:0] out_data;

assign out_data = 
				(in_data == 7'd00) ?  14'd07540 : 
				(in_data == 7'd01) ?  14'd07110 : 
				(in_data == 7'd02) ?  14'd06704 : 
				(in_data == 7'd03) ?  14'd06321 : 
				(in_data == 7'd04) ?  14'd05959 : 
				(in_data == 7'd05) ?  14'd05619 : 
				(in_data == 7'd06) ?  14'd05298 : 
				(in_data == 7'd07) ?  14'd04995 : 
				(in_data == 7'd08) ?  14'd04710 : 
				(in_data == 7'd09) ?  14'd04441 : 
				(in_data == 7'd010) ?  14'd04187 : 
				(in_data == 7'd011) ?  14'd03948 : 
				(in_data == 7'd012) ?  14'd03722 : 
				(in_data == 7'd013) ?  14'd03510 : 
				(in_data == 7'd014) ?  14'd03309 : 
				(in_data == 7'd015) ?  14'd03120 : 
				(in_data == 7'd016) ?  14'd02942 : 
				(in_data == 7'd017) ?  14'd02774 : 
				(in_data == 7'd018) ?  14'd02615 : 
				(in_data == 7'd019) ?  14'd02466 : 
				(in_data == 7'd020) ?  14'd02325 : 
				(in_data == 7'd021) ?  14'd02192 : 
				(in_data == 7'd022) ?  14'd02067 : 
				(in_data == 7'd023) ?  14'd01949 : 
				(in_data == 7'd024) ?  14'd01838 : 
				(in_data == 7'd025) ?  14'd01733 : 
				(in_data == 7'd026) ?  14'd01634 : 
				(in_data == 7'd027) ?  14'd01540 : 
				(in_data == 7'd028) ?  14'd01452 : 
				(in_data == 7'd029) ?  14'd01369 : 
				(in_data == 7'd030) ?  14'd01291 : 
				(in_data == 7'd031) ?  14'd01217 : 
				(in_data == 7'd032) ?  14'd01148 : 
				(in_data == 7'd033) ?  14'd01082 : 
				(in_data == 7'd034) ?  14'd01020 : 
				(in_data == 7'd035) ?  14'd0962 : 
				(in_data == 7'd036) ?  14'd0907 : 
				(in_data == 7'd037) ?  14'd0855 : 
				(in_data == 7'd038) ?  14'd0807 : 
				(in_data == 7'd039) ?  14'd0760 : 
				(in_data == 7'd040) ?  14'd0717 : 
				(in_data == 7'd041) ?  14'd0676 : 
				(in_data == 7'd042) ?  14'd0637 : 
				(in_data == 7'd043) ?  14'd0601 : 
				(in_data == 7'd044) ?  14'd0567 : 
				(in_data == 7'd045) ?  14'd0534 : 
				(in_data == 7'd046) ?  14'd0504 : 
				(in_data == 7'd047) ?  14'd0475 : 
				(in_data == 7'd048) ?  14'd0448 : 
				(in_data == 7'd049) ?  14'd0422 : 
				(in_data == 7'd050) ?  14'd0398 : 
				(in_data == 7'd051) ?  14'd0375 : 
				(in_data == 7'd052) ?  14'd0354 : 
				(in_data == 7'd053) ?  14'd0334 : 
				(in_data == 7'd054) ?  14'd0315 : 
				(in_data == 7'd055) ?  14'd0297 : 
				(in_data == 7'd056) ?  14'd0280 : 
				(in_data == 7'd057) ?  14'd0264 : 
				(in_data == 7'd058) ?  14'd0249 : 
				(in_data == 7'd059) ?  14'd0234 : 
				(in_data == 7'd060) ?  14'd0221 : 
				(in_data == 7'd061) ?  14'd0208 : 
				(in_data == 7'd062) ?  14'd0197 : 
				(in_data == 7'd063) ?  14'd0185 : 
				(in_data == 7'd064) ?  14'd0175 : 
				(in_data == 7'd065) ?  14'd0165 : 
				(in_data == 7'd066) ?  14'd0155 : 
				(in_data == 7'd067) ?  14'd0146 : 
				(in_data == 7'd068) ?  14'd0138 : 
				(in_data == 7'd069) ?  14'd0130 : 
				(in_data == 7'd070) ?  14'd0123 : 
				(in_data == 7'd071) ?  14'd0116 : 
				(in_data == 7'd072) ?  14'd0109 : 
				(in_data == 7'd073) ?  14'd0103 : 
				(in_data == 7'd074) ?  14'd097 : 
				(in_data == 7'd075) ?  14'd091 : 
				(in_data == 7'd076) ?  14'd086 : 
				(in_data == 7'd077) ?  14'd081 : 
				(in_data == 7'd078) ?  14'd077 : 
				(in_data == 7'd079) ?  14'd072 : 
				(in_data == 7'd080) ?  14'd068 : 
				(in_data == 7'd081) ?  14'd064 : 
				(in_data == 7'd082) ?  14'd061 : 
				(in_data == 7'd083) ?  14'd057 : 
				(in_data == 7'd084) ?  14'd054 : 
				(in_data == 7'd085) ?  14'd051 : 
				(in_data == 7'd086) ?  14'd048 : 
				(in_data == 7'd087) ?  14'd045 : 
				(in_data == 7'd088) ?  14'd043 : 
				(in_data == 7'd089) ?  14'd040 : 
				(in_data == 7'd090) ?  14'd038 : 
				(in_data == 7'd091) ?  14'd036 : 
				(in_data == 7'd092) ?  14'd034 : 
				(in_data == 7'd093) ?  14'd032 : 
				(in_data == 7'd094) ?  14'd030 : 
				(in_data == 7'd095) ?  14'd028 : 
				(in_data == 7'd096) ?  14'd027 : 
				(in_data == 7'd097) ?  14'd025 : 
				(in_data == 7'd098) ?  14'd024 : 
				(in_data == 7'd099) ?  14'd022 : 
				(in_data == 7'd0100) ?  14'd021 : 
				(in_data == 7'd0101) ?  14'd020 : 
				(in_data == 7'd0102) ?  14'd019 : 
				(in_data == 7'd0103) ?  14'd018 : 
				(in_data == 7'd0104) ?  14'd017 : 
				(in_data == 7'd0105) ?  14'd016 : 
				(in_data == 7'd0106) ?  14'd015 : 
				(in_data == 7'd0107) ?  14'd014 : 
				(in_data == 7'd0108) ?  14'd013 : 
				(in_data == 7'd0109) ?  14'd012 : 
				(in_data == 7'd0110) ?  14'd012 : 
				(in_data == 7'd0111) ?  14'd011 : 
				(in_data == 7'd0112) ?  14'd010 : 
				(in_data == 7'd0113) ?  14'd010 : 
				(in_data == 7'd0114) ?  14'd09 : 
				(in_data == 7'd0115) ?  14'd09 : 
				(in_data == 7'd0116) ?  14'd08 : 
				(in_data == 7'd0117) ?  14'd08 : 
				(in_data == 7'd0118) ?  14'd07 : 
				(in_data == 7'd0119) ?  14'd07 : 
				(in_data == 7'd0120) ?  14'd06 : 
				(in_data == 7'd0121) ?  14'd06 : 
				(in_data == 7'd0122) ?  14'd06 : 
				(in_data == 7'd0123) ?  14'd05 : 
				(in_data == 7'd0124) ?  14'd05 : 
				(in_data == 7'd0125) ?  14'd05 : 
				(in_data == 7'd0126) ?  14'd05 : 
				(in_data == 7'd0127) ?  14'd04 : 15'd0 ;
									 
endmodule